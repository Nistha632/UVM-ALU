interface alu_interface;
  
  logic [2 : 0 ]  mode;
  logic [3 : 0 ]   a,b;
  logic [7 : 0 ]     y;
 
endinterface


